interface AES_intf();
import shared_pkg::*;
    logic [127:0] in;
    logic [127:0] key;
    logic [127:0] out;
endinterface //AES