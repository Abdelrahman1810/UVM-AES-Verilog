package shared_pkg;
parameter N=128;
parameter Nr=10;
parameter Nk=4;
parameter LOOP = 100;
endpackage